module UART_RX #(parameter CLKS_PER_BIT = 5200)(
  input        i_rx_data,
  input        i_clock,
  output       o_rx_dv,
  output [7:0] o_rx_data);
  
  parameter S_IDLE      = 3'b000;
  parameter S_START_BIT = 3'b001;
  parameter S_DATA_BITS = 3'b010;
  parameter S_STOP_BIT  = 3'b011;
  parameter S_CLEANUP   = 3'b100;
  
  reg [7:0] r_byte;
  reg [7:0] clk_count;
  reg [2:0] bit_index;
  reg [2:0] state;
  reg       r_rx_dv;
  reg       r_data;
  reg       r_data_r;
  
  always@(posedge i_clock)		// we are using dual flip flops to avoid metastability
    begin
      r_data_r <= i_rx_data;
      r_data   <= r_data_r;
    end
  
  
  always@(posedge i_clock)
    begin
      case(state)
        
        S_IDLE :
          begin
            clk_count <= 0;
            bit_index <= 0;
            r_rx_dv   <= 1'b0;
            
            if(i_rx_data == 1'b0)		// start bit detection
              state    <= S_START_BIT;
            else
              state <= S_IDLE;
          end
        
        S_START_BIT :
          begin
            if(clk_count == (CLKS_PER_BIT - 1)/2)	// finding the middle of start bit
              begin
                if(r_data == 1'b0)
                  begin
                    clk_count <= 0;				// resetting counter
                    state     <= S_DATA_BITS;
                  end
                else
                  begin
                    state  <= S_IDLE;
                  end
              end
            else
              begin
                clk_count <= clk_count + 1;
                state     <= S_START_BIT;
              end
          end
        
        S_DATA_BITS :
          begin
            if(clk_count < CLKS_PER_BIT - 1)
              begin
                clk_count <= clk_count + 1;
                state     <= S_DATA_BITS;
              end
            else
              begin
                clk_count         <= 0;
                r_byte[bit_index] <= r_data;
                
                if(bit_index < 7)
                  begin
                    bit_index <= bit_index + 1;
                    state     <= S_DATA_BITS;
                  end
                else
                  begin
                    bit_index <= 0;
                    state     <= S_STOP_BIT;
                  end
              end
          end
        
        S_STOP_BIT :
          begin
            if(clk_count < CLKS_PER_BIT - 1)
              begin
                clk_count <= clk_count + 1;
                state     <= S_STOP_BIT;
              end
            else
              begin
                clk_count <= 0;
                r_rx_dv   <= 1'b1;
                state     <= S_CLEANUP;
              end
          end
        
        S_CLEANUP :
          begin
            r_rx_dv <= 1'b0;
            state   <= S_IDLE;
          end
        
        default :
          state <= S_IDLE;
      endcase
    end
  
  assign o_rx_dv   = r_rx_dv;
  assign o_rx_data = r_byte;
  
endmodule
